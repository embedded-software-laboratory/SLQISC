module vgabox
#(
    parameter SYMBOLS = 4,
	 parameter TOP = 0,
	 parameter LEFT = 0
)
(
  input [8:0] curRow,
  input [9:0] curCol,
  input [7*SYMBOLS-1:0] characters,
  output pixel
);


wire [8:0] charRow;
wire [9:0] charCol;
	
wire [8:0] inCharRow;
wire [9:0] inCharCol;
	
wire [49:0] pixelGrid;
wire [7:0] pixelRow;
wire superpixel;
wire outbox;

assign charCol = (curCol - (LEFT-8)) >> 5;
assign inCharCol = ((curCol - (LEFT-8)) & 9'h1f) >> 2;
assign inCharRow = (curRow - TOP) >> 2;
assign pixelGrid = {charMap(characters[charCol * 7 +: 7]), 5'b0};
assign pixelRow = {pixelGrid[inCharRow*5 +: 5], 3'b0};
assign superpixel = pixelRow[inCharCol] && TOP + 4 <= curRow && curRow < TOP + 40 && LEFT + 4 <= curCol && curCol < LEFT + 32*SYMBOLS-8;
assign outbox = TOP <= curRow && curRow < TOP+44 && LEFT <= curCol && curCol < LEFT+32*SYMBOLS-4;
assign pixel = !superpixel && outbox;

//" ABCDEFGHIJKLMNOPQRSTUVWXYZ!0123456789abcdefghijklmnopqrstuvwxyz+-"
function [44:0] charMap (input[6:0] chr);
  begin
  case(chr)
    00: charMap=45'b0;
	 01: charMap=45'b10001_10001_10001_10001_11111_10001_10001_10001_11111;
	 02: charMap=45'b01111_10001_10001_10001_01111_10001_10001_10001_01111;
	 03: charMap=45'b11110_00001_00001_00001_00001_00001_00001_00001_11110;
	 04: charMap=45'b01111_10001_10001_10001_10001_10001_10001_10001_01111;
	 05: charMap=45'b11111_00001_00001_00001_00111_00001_00001_00001_11111;
	 06: charMap=45'b00001_00001_00001_00001_00111_00001_00001_00001_11111;
	 07: charMap=45'b01110_10001_10001_10001_01101_00001_10001_10001_01110;
	 08: charMap=45'b10001_10001_10001_10001_11111_10001_10001_10001_10001;
	 09: charMap=45'b00100_00100_00100_00100_00100_00100_00100_00100_00100;
	 12: charMap=45'b11111_00001_00001_00001_00001_00001_00001_00001_00001;
	 14: charMap=45'b10001_11001_11001_10101_10101_10101_10011_10011_10001;
	 15: charMap=45'b01110_10001_10001_10001_10001_10001_10001_10001_01110;
	 18: charMap=45'b10001_01001_00101_00011_01111_10001_10001_10001_01111;
	 19: charMap=45'b01110_10001_10000_01000_00100_00010_00001_10001_01110;
	 20: charMap=45'b00100_00100_00100_00100_00100_00100_00100_00100_11111;
	 21: charMap=45'b01110_10001_10001_10001_10001_10001_10001_10001_10001;
	 22: charMap=45'b00100_01010_10001_10001_10001_10001_10001_10001_10001;
	 23: charMap=45'b10001_11011_10101_10101_10101_10001_10001_10001_10001;
	 25: charMap=45'b00100_00100_00100_00100_00100_01010_01010_10001_10001;
	 27: charMap=45'b00100_00000_00000_00100_00100_00100_00100_00100_00100;
	 28: charMap=45'b01110_10001_10001_10101_10101_10101_10001_10001_01110;
	 29: charMap=45'b10000_10000_10000_10000_10001_10010_10100_11000_10000;
	 30: charMap=45'b11111_00010_00100_01000_10000_10001_10001_10001_01110;
	 31: charMap=45'b01110_10001_10000_10000_01110_10000_10000_10001_01110;
	 32: charMap=45'b00100_00100_00100_00100_11111_00101_00101_00101_00101;
	 33: charMap=45'b01110_10001_10000_10000_01111_00001_00001_00001_11111;
	 34: charMap=45'b01110_10001_10001_10001_01111_00001_00001_00001_01110;
	 35: charMap=45'b00100_00100_00100_00100_00100_01000_01000_10000_11111;
	 36: charMap=45'b01110_10001_10001_10001_01110_10001_10001_10001_01110;
	 37: charMap=45'b01110_10001_10000_10000_11110_10001_10001_10001_01110;
    default: charMap=45'b11111_11111_11111_11111_11111_11111_11111_11111_11111;
  endcase
  end
endfunction


endmodule